DIFF���E    �DM�/	1b�ID;�d�� d�  � �n�  `�+����^�ľN�G桎4*�bĊi.s�x�<��zW@@*�*+��U���ђ5�i��^m���{#җ5�&�;5�B���#�7H���bLL���v�-�8�Q=ѥ5R�JGC�\S�	^��:Ŏ�[�p���T%j�*��y��f$���n�ϕY���Dʕ���fS(~@�Z䦦02)_yP���\�E�;�|�*���O��Q8ba�/OC�V��fRX��v�Y��[��ڭ��R+t�[ B��S=�)d	;��*lߵ;�Ľ.U;��⾖%	��z�VVNm���W<�O���wKK�rr2� ���H���;��n���p�| ����#%�~�\���xb�A�S~������6/}�7�.��Lm�"]h{Y��4{�n��TT�#��}!��8�����+��'QL~��۬��uC�l��l�Y�>��%,�ф�I�P�E��p�	�"��P*�inp��M���\�ǒ��8�m�Kd� ƥ��w%?���kc��yGyX�[��9��z����3G)E��m�S� 